module vga_pic(
	vga_clk				,
	rst_n				,
	pix_x				,
	pix_y				,

	pix_data			 
);
	input		 		vga_clk			;			
	input		 		rst_n			;			
	input  [9:0] 		pix_x			;			
	input  [9:0] 		pix_y			;			
	output [15:0]		pix_data		;

	reg    [15:0]		pix_data		;

	parameter			CHAR_B_H 		= 10'd192,
						CHAR_B_V		= 10'd208;

	parameter			CHAR_W			= 10'd256,
						CHAR_H			= 10'd64 ;
	parameter			BLACK			= 16'h0000,
						GOLDEN			= 16'hFEC0;
	

	reg   [255:0]		char	[63:0]	;
	wire  [9:0]			char_x			;
	wire  [9:0]			char_y			;

	assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
					&& ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H)))) ? (pix_x - CHAR_B_H) : 10'h3ff;
	assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W))) && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H)))) ? (pix_y - CHAR_B_V) : 10'h3ff;

	always@(posedge vga_clk)
	begin
		char[00]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[01]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[02]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[03]	<= 256'h000000700000000000000000000000000000000300000000000000007C000000;
		char[04]	<= 256'h0000003E0000000000000000000000000000200380000000000010003F000000;
		char[05]	<= 256'h0000003E00000000000000007800000000003803E000000000001C001F800000;
		char[06]	<= 256'h0000003C000000000000000FFC00000000003C03C000000000003E000FC00000;
		char[07]	<= 256'h0000001C00000000000011FF7F000000000078078000000000003E0403C00000;
		char[08]	<= 256'h0000001C1E00000000001F803F00000000007007800000000000780F00C00000;
		char[09]	<= 256'h0000001C0F80000000001E001E0000000000F00F000000000000F00F80000000;
		char[10]	<= 256'h0000001C07C0000000000E001E0000000000E00E007000000001C00F00000000;
		char[11]	<= 256'h0000000C03E0000000000E003C0000000001C01C03FC00000007021E00000000;
		char[12]	<= 256'h0000000C03E0000000000F0F3C0000000001C01CFFFE0000000E07FC00000000;
		char[13]	<= 256'h0000000C00C00000000007FF380000000003803FE03F0000001801F800000000;
		char[14]	<= 256'h0000070E00000000000007F83800000000070070003F00000000007C00000000;
		char[15]	<= 256'h00000F8E000000000000070038000000000780E000780000000000FF00000000;
		char[16]	<= 256'h00001F86000000000000030038000000000F80C180600000000001E7C0000000;
		char[17]	<= 256'h00003E06000000000000030030000000001DC180F0C00000000003C1F0000000;
		char[18]	<= 256'h000078060000000000000300300000000038C300E000000000000700FE000000;
		char[19]	<= 256'h0000E007000000000000030FF00000000070C400E000000000000E303FC00000;
		char[20]	<= 256'h0003F0070F000000000003FFE00000000060C0006000000000001C3C0FFC0000;
		char[21]	<= 256'h000038037F000000000001C00000000000C0C040630000000000787C07FFF000;
		char[22]	<= 256'h00003C07FC0000000000010001E000000180C04061F000000000F07FC1FFF800;
		char[23]	<= 256'h00001C3FE0000000000000001FF000000200C0C060FC00000001C0F7E07F0000;
		char[24]	<= 256'h00001DFF8000000000000001FFF800000000C1C0607C0000000781C3F0000000;
		char[25]	<= 256'h00001FF1808000000000003FFFE000000001C1C0603E0000001E0783E0000000;
		char[26]	<= 256'h00007F81C0E00000000007FF000000000001C3C0601E000000780F0780000000;
		char[27]	<= 256'h0007FC01C0F000000000FFFE000000000001C380F00E000001E01E0F00000000;
		char[28]	<= 256'h00FFCC00C0F0000000FFFE0E000000000001C180F000000006007B9E00000000;
		char[29]	<= 256'h007E0C00E1E0000000FFC00E000000000003C00FF00000000001C3FC00000000;
		char[30]	<= 256'h00100C6061E00000003E200E0000000000038007E0000000000001F800000000;
		char[31]	<= 256'h00000D8063C000000000780E0C00000000038001E0000000000001E700000000;
		char[32]	<= 256'h00000F00738000000000780E7F00000000018001E0000000000003C780000000;
		char[33]	<= 256'h00001E00370000000000780FFF00000000018000C07E000000000F8F80000000;
		char[34]	<= 256'h0000FC003F0000000000F80FF800000000000070403FC00000003E1FFE000000;
		char[35]	<= 256'h0003FC001E0000000001F80E000000000008007C001FE0000000783CFF000000;
		char[36]	<= 256'h001F9C003C0000000001FC0E000000000008003E0007F0000001E0781F800000;
		char[37]	<= 256'h00FE1C003E0000000003C70E000000000008001F0003F000000780F01E000000;
		char[38]	<= 256'h07F81C007F0000000007838E000000000018200F0000F000001803E03C000000;
		char[39]	<= 256'h07F01C01E7000000000701EC0000000000183003000078000000078078000000;
		char[40]	<= 256'h01C01C03C7800000000F00FC00000000001810000200000000001EC0F0000000;
		char[41]	<= 256'h00001C0F03C02000001E003C000000000038180001000000000078E1E0000000;
		char[42]	<= 256'h00001C1C01E02000003C001F0000000000780C00018000000001C073C0000000;
		char[43]	<= 256'h00001C6000F020000078000FC000000000780E0000C000000000007780000000;
		char[44]	<= 256'h0003FC000078200000E00003F000000000F8078000E000000000003F00000000;
		char[45]	<= 256'h0001F800007C600001C00001FF00000000F003E000F800000000003C00000000;
		char[46]	<= 256'h0000F800003FF00007800000FFF80000006001FFC7FC0000000000F800000000;
		char[47]	<= 256'h00007800001FF0000E0000007FFFF000004000FFFFFC0000000003E000000000;
		char[48]	<= 256'h000030000007F000000000001FFFFC000000003FFFF8000000000FC000000000;
		char[49]	<= 256'h000020000003F000000000000FFFC00000000007FF80000000003F0000000000;
		char[50]	<= 256'h000000000001F0000000000003FC000000000000000000000000FC0000000000;
		char[51]	<= 256'h0000000000007000000000000000000000000000000000000007E00000000000;
		char[52]	<= 256'h000000000000000000000000000000000000000000000000007F000000000000;
		char[53]	<= 256'h0000000000000000000000000000000000000000000000000080000000000000;
		char[54]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[55]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[56]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[57]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[58]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[59]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[60]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[61]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[62]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[63]	<= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	end

	always  @(posedge vga_clk or negedge rst_n)begin
		if(rst_n==1'b0)begin
			pix_data	<= BLACK;
		end
		else if(((pix_x >= CHAR_B_H - 1'b1) && (pix_x < (CHAR_B_H + CHAR_W - 1'b1)))
					&& ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H)))
					&& (char[char_y][10'd255 - char_x] == 1'b1))begin
			pix_data	<= GOLDEN;
		end
		else begin
			pix_data	<= BLACK;
		end
	end

endmodule

