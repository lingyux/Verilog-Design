library verilog;
use verilog.vl_types.all;
entity ring_tb is
end ring_tb;
