library verilog;
use verilog.vl_types.all;
entity tb_my_vga is
end tb_my_vga;
