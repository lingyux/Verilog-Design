library verilog;
use verilog.vl_types.all;
entity divider_tb is
end divider_tb;
