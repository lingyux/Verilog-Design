library verilog;
use verilog.vl_types.all;
entity Rs232_tb is
end Rs232_tb;
