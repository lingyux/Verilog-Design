library verilog;
use verilog.vl_types.all;
entity tb_tft_colorbar is
end tb_tft_colorbar;
