library verilog;
use verilog.vl_types.all;
entity tb_led_ctrl is
end tb_led_ctrl;
